library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity top_module is
  port (
    clk          : in  std_logic;
    reset_n      : in  std_logic;
    rx           : in  std_logic;
    tx           : out std_logic
  );
end top_module;

architecture rtl of top_module is

  -- Sinais internos
  signal baud_tick     : std_logic;

  -- Interface UART RX -> FIFO TX
  signal s_axis_tdata  : std_logic_vector(7 downto 0);
  signal s_axis_tvalid : std_logic;
  signal s_axis_tready : std_logic;

  -- FIFO TX -> FIFO RX
  signal fifo_tdata0    : std_logic_vector(7 downto 0);
  signal fifo_tvalid0   : std_logic;
  signal fifo_tready0   : std_logic;

  -- FIFO RX -> UART TX
  signal fifo_tdata1    : std_logic_vector(7 downto 0);
  signal fifo_tvalid1   : std_logic;
  signal fifo_tready1   : std_logic;

  -- Controle do UART TX
  signal tx_busy        : std_logic;
  signal tx_start       : std_logic;

  -- Sinais "Dummy" (para conectar as saídas de debug)
  signal ignore_data    : std_logic_vector(7 downto 0);
  signal ignore_valid   : std_logic;
  signal ignore_ready   : std_logic;
  signal ignore_error1  : std_logic;
  signal ignore_error2  : std_logic;
  signal ignore_busy    : std_logic;

  -- NOVOS SINAIS para conectar o Filtro
  signal filter_out_data  : std_logic_vector(7 downto 0);
  signal filter_out_valid : std_logic;
  signal filter_out_ready : std_logic;

begin

  -- 1. Gerador de Baud Rate (Lembre-se: 25MHz para Colorlight i9+)
  baud_gen_inst : entity work.baud_gen
    generic map (
      CLK_FREQ  => 25_000_000, 
      BAUD_RATE => 115200      
    )
    port map (
      clk       => clk,
      reset_n   => reset_n,
      baud_tick => baud_tick
    );

  -- -- 2. Receptor UART
  -- uart_rx_inst : entity work.uart_rx
  --   generic map (
  --     DATA_BITS => 8,
  --     STOP_BITS => 1,
  --     PARITY    => "NONE"
  --   )
  --   port map (
  --     clk          => clk,
  --     reset_n      => reset_n,
  --     rx           => rx,
  --     baud_tick    => baud_tick,
  --     axis_tdata   => s_axis_tdata,
  --     axis_tvalid  => s_axis_tvalid,
  --     axis_tready  => s_axis_tready,
  --     -- Conectamos em sinais internos que não vão a lugar nenhum
  --     frame_error  => ignore_error1,
  --     parity_error => ignore_error2,
  --     busy         => ignore_busy
  --   );

  -- 2. Receptor UART (Atualizado com timer interno)
  uart_rx_inst : entity work.uart_rx
    generic map (
      DATA_BITS => 8,
      STOP_BITS => 1,
      PARITY    => "NONE",
      CLK_FREQ  => 25_000_000, -- Configure para o clock da Colorlight i9+
      BAUD_RATE => 115_200
    )
    port map (
      clk          => clk,
      reset_n      => reset_n,
      rx           => rx,
      -- baud_tick => baud_tick, -- REMOVIDO: RX gera seu proprio timing
      axis_tdata   => s_axis_tdata,
      axis_tvalid  => s_axis_tvalid,
      axis_tready  => s_axis_tready,
      frame_error  => ignore_error1,
      parity_error => ignore_error2,
      busy         => ignore_busy
    );

  -- 3. FIFO RX (TX do lado da FPGA, RX do lado da UART)
  fifo_rx_inst : entity work.fifo_UART
    generic map ( DATA_WIDTH => 8, DEPTH => 4096 ) -- Mantendo o buffer grande!
    port map (
      clk          => clk,
      reset_n      => reset_n,
      axis_tdata   => s_axis_tdata,
      axis_tvalid  => s_axis_tvalid,
      axis_tready  => s_axis_tready,
      -- A SAÍDA DA FIFO AGORA VAI PARA O FILTRO
      fifo_tdata   => fifo_tdata0,
      fifo_tvalid  => fifo_tvalid0,
      fifo_tready  => fifo_tready0 
    );

  -- 3.5 NOVO BLOCO: FILTRO DE IMAGEM
  img_filter_inst : entity work.image_filter
    generic map (
      IMG_WIDTH  => 150 -- Tem que bater com o Python
    )
    port map (
      -- (sinais continuam iguais)
      clk           => clk,
      reset_n       => reset_n,
      s_axis_tdata  => fifo_tdata0,
      s_axis_tvalid => fifo_tvalid0,
      s_axis_tready => fifo_tready0,
      m_axis_tdata  => filter_out_data,
      m_axis_tvalid => filter_out_valid,
      m_axis_tready => filter_out_ready
    );

  -- 4. FIFO TX (Buffer para saída)
  fifo_tx_inst : entity work.fifo_UART
    generic map ( DATA_WIDTH => 8, DEPTH => 4096 )
    port map (
      clk          => clk,
      reset_n      => reset_n,
      -- A ENTRADA VEM DO FILTRO
      axis_tdata   => filter_out_data,
      axis_tvalid  => filter_out_valid,
      axis_tready  => filter_out_ready,
      
      fifo_tdata   => fifo_tdata1,
      fifo_tvalid  => fifo_tvalid1,
      fifo_tready  => fifo_tready1
    );

  -- -- 3. FIFO Intermediária 1 (TX)
  -- fifo_rx_inst : entity work.fifo_UART
  --   generic map ( DATA_WIDTH => 8, DEPTH => 4096 )
  --   port map (
  --     clk          => clk,
  --     reset_n      => reset_n,
  --     axis_tdata   => s_axis_tdata,
  --     axis_tvalid  => s_axis_tvalid,
  --     axis_tready  => s_axis_tready,
  --     fifo_tdata   => fifo_tdata0,
  --     fifo_tvalid  => fifo_tvalid0,
  --     fifo_tready  => fifo_tready0
  --   );

  -- -- 4. FIFO Intermediária 2 (RX)
  -- fifo_tx_inst : entity work.fifo_UART
  --   generic map ( DATA_WIDTH => 8, DEPTH => 4096 )
  --   port map (
  --     clk          => clk,
  --     reset_n      => reset_n,
  --     axis_tdata   => fifo_tdata0,
  --     axis_tvalid  => fifo_tvalid0,
  --     axis_tready  => fifo_tready0,
  --     fifo_tdata   => fifo_tdata1,
  --     fifo_tvalid  => fifo_tvalid1,
  --     fifo_tready  => fifo_tready1
  --   );

  -- 5. Lógica de Controle
  process(fifo_tvalid1, tx_busy)
  begin
    if (fifo_tvalid1 = '1' and tx_busy = '0') then
      tx_start     <= '1';
      fifo_tready1 <= '1';
    else
      tx_start     <= '0';
      fifo_tready1 <= '0';
    end if;
  end process;

  -- 6. Transmissor UART
  uart_tx_inst : entity work.uart_tx
    generic map (
      DATA_BITS => 8,
      STOP_BITS => 1,
      PARITY    => "NONE"
    )
    port map (
      clk       => clk,
      reset_n   => reset_n,
      baud_tick => baud_tick,
      tx_start  => tx_start,
      tx_data   => fifo_tdata1,
      tx        => tx,
      busy      => tx_busy
    );

end rtl;