module top (
  input sys_clk
);
  
endmodule