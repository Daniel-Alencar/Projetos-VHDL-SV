module pll(
  input sys_clk,
  output pll_clk, pll_lock
);
endmodule