library ieee;
use ieee.std_logic_1164.all;

package types_pkg is
    type int_array is array (natural range <>) of integer;
end package;
